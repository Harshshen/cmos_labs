** Y = (AB + C(D + E))'
.subckt pass_and 1 2 3 4
.model nmod nmos level = 54 version = 4.7
M1 2 3 4 4 nmod w = 100u l = 10u
M2 1 2 4 4 nmod w = 100u l = 10u
.ends
.subckt pass_or 1 2 3 4
.model nmod nmos level = 54 version = 4.7
M1 2 2 4 4 nmod w = 100u l = 10u
M2 1 3 4 4 nmod w = 100u l = 10u
.ends
.subckt pass_inverter 1 2 3
.model nmod nmos level = 54 version = 4.7
.model pmod pmos level = 54 version = 4.7
M1 3 1 2 2 pmod w = 100u l = 10u
M2 3 1 0 0 nmod w = 100u l = 10u
.ends
Va 11 0 pulse(0 5 0 0 0 10m 20m)
Vb 12 0 dc 5V
Vc 13 0 dc 5V
Vd 14 0 dc 5V
Ve 15 0 dc 5V
Vdd 2 0 dc 5V
Xb 12 2 20 pass_inverter
Xc 13 2 16 pass_inverter
Xe 15 2 17 pass_inverter
Xcanddore 19 2 22 pass_inverter
Xaandb 11 12 20 21 pass_and
Xdore 14 15 17 18 pass_or
Xdoreandc 18 13 16 19 pass_and
Xaandbordore 21 19 22 23 pass_or
.tran 0.1m 500m
.control
run
plot V(11) V(12) V(13) V(14) V(15) V(23)
.endc
.end
