* 2 input and gate*
vd 5 0 dc 5v
va 3 0 dc 5v
vb 1 0 pulse(0 5 0 0 0 5m 10m)

.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
M1 4 3 2 0 nmod w=100u l=10u
M2 2 3 0 0 nmod w=100u l=10u
M3 4 1 5 0 pmod w=100u l=10u
M4 4 1 5 0 pmod w=100u l=10u

.tran 0.1m 80m
.control
run
plot V(1) V(4)
.endc
.end
