*MUX USING TRANSMISSION GATE*
.subckt inverter 1 2 3
M1 3 1 0 0 nmod w=100u l=10u
M2 3 1 2 2 pmod w=100u l=10u
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
.ends
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
Va 10 0 dc 5
Vb 11 0 dc 0
Vd1 2 0 dc 5
xs 3 2 4 inverter
Vs 3 0 pulse (0 5 0 0 0 10m 20m)
M1 1 4 5 5 nmod w=100u l=10u
M2 1 3 5 5 pmod w=100u l=10u
M3 2 3 5 5 nmod w=100u l=10u
M4 2 4 5 5 pmod w=100u l=10u
.tran 0.1m 40m
.control
run
plot V(3) V(5)
.endc
.end